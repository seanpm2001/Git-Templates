// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 1
// For: /SNU/2D/ProgrammingTools/IDE/Verilog-AMS/
// About:
// -- I decided to make Verilog-AMS the main project language file for this project (SNU / 2D / Programming Tools / IDE / Grammatical-Framework) as this is a Verilog-AMS IDE, and it needs its main language to be represented here.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 01'00000000 // Random data to test syntax
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: Verilog-AMS source file (*.v *.vh)
// File version: 1 (2022, Tuesday, October 25th at 12:58 pm PST)
// Line count (including blank lines and compiler line): 16
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script
