-- Start of script

-- I have chosen VHDL as the 3rd project language file for this project (Seanpm2001/OuterVM-Mouse) as along with Assembly, it is needed for hardware virtualization.

-- File info

-- File version: 1 (Sunday, 2021 October 24th at 5:29 pm)
-- File type: Virtual Hard Disk Language (VHDL) Source file (*.vhdl, *.vhd, *.vdi)
-- Line count (including blank lines and compiler line): 12

-- End of script
