-- Start of script
-- This project (RecursionBot) contains source code in Virtual Hard Disk Language (VHDL) format, as it is one of the 9 languages needed to be used to build the program.");
-- File version: 1 (Wednesday, March 3rd 2021 at 6:54 pm)
-- File type: Virtual Hard Disk Language (VHDL) Source file (*.vhdl)
-- Line count (including blank lines and compiler line): 7
-- End of script
