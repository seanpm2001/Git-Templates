-- Start of script

-- I decided to make VHDL the main project language file for this project (Seanpm2001/Learn-VHDL) as VHDL is the language this project is dedicated to, because this project is about learning the VHDL programming language. It only makes sense to make VHDL the official language for this project.

-- File info

-- File version: 1 (Friday, 2021 November 26th at 6:28 pm)
-- File type: Virtual Hard Disk Language (VHDL) Source file (*.vhdl, *.vhd, *.vdi)
-- Line count (including blank lines and compiler line): 12

-- End of script

