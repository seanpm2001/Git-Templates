// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 1
// For: Metro Techno
// I decided to make Verilog the first project language file for this project (Seanpm2001/MetroTechno) as Verilog is the primary language used for system programming throughout the Metro Techno system map. Although 7 other languages are planned to be used, Verilog comes first. It is getting its own project language file, starting here.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 01'00000000 // Random data to test syntax (also: 0 in binary)
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: Verilog source file (*.v *.vh)
// File version: 1 (2022, Wednesday, September 7th at 7:10 pm PST)
// Line count (including blank lines and compiler line): 15
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script
