// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 4
// For: BootDown
// I have decided to make SystemVerilog the 4th project language file for this project (BootDown) as it is a good alternative scripting language for the low-level parts of the system this project is designed for. It is also a newer version of Verilog that I also want to use.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 4'00000100 // Random data to test syntax
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: SystemVerilog source file (*.sv *.svh)
// File version: 1 (Monday, 2021 September 20th at 2:16 pm)
// Line count (including blank lines and compiler line): 15
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script

