-- Start of script

-- Notes
-- I don't know how to make strings in VHDL, so comments will do for now

-- Project language file 1
-- For: /SNU/2D/ProgrammingTools/IDE/VHDL/
-- About:
-- I decided to make VHDL the main project language file for this project (SNU / 2D / Programming Tools / IDE / VHDL) as this is a VHDL IDE, and it needs its main language to be represented here.

-- File info

-- File version: 1 (2022, Sunday, October 16th at 5:32 pm PST)
-- File type: Virtual Hard Disk Language (VHDL) Source file (*.vhdl, *.vhd, *.vdi)
-- Line count (including blank lines and compiler line): 18

-- End of script
