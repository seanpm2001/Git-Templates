// Start of script */

// Project language file 1
// For: /SNU/2D/ProgrammingTools/IDE/Verilog/
// About:
// I decided to make Verilog the main project language file for this project (SNU / 2D / Programming Tools / IDE / Verilog) as this is a Verilog IDE, and it needs its main language to be represented here.

module main;
  initial
    begin
      $display("Project language file 1");
      $display("For: /SNU/2D/ProgrammingTools/IDE/Verilog/");
      $display("About:");
      $display("I decided to make Verilog the main project language file for this project (SNU / 2D / Programming Tools / IDE / Verilog) as this is a Verilog IDE, and it needs its main language to be represented here.");
      $finish;
    end
endmodule

// File info
// File type: Verilog source file (*.v *.vh)
// File version: 1 (2022, Saturday, November 5th at 11:01 pm PST)
// Line count (including blank lines and compiler line): 25

// End of script */
