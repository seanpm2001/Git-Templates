-- Start of script
-- I have chosen VHDL as the 2nd project language file for this project (BootDown) as along with Assembly, it is needed for hardware virtualization.
-- File version: 1 (Monday, 2021 September 20th at 1:59 pm)
-- File type: Virtual Hard Disk Language (VHDL) Source file (*.vhdl, *.vhd, *.vdi)
-- Line count (including blank lines and compiler line): 7
-- End of script
