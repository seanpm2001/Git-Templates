// Start of script */

// Project language file 1
// For: seanpm2001/Learn-Verilog-AMS
// About:
// I decided to make Verilog-AMS the main project language file for this project (Seanpm2001/Learn-Verilog-AMS) as Verilog-AMS is the language this project is dedicated to, because this project is about learning the Verilog-AMS programming language. It only makes sense to Verilog-AMS the official language for this project. It is getting its own project language file, starting here.

module main;
  initial
    begin
      $display("Project language file 1");
      $display("For: seanpm2001/Learn-Verilog-AMS");
      $display("About:");
      $display("I decided to make Verilog-AMS the main project language file for this project (Seanpm2001/Learn-Verilog-AMS) as Verilog-AMS is the language this project is dedicated to, because this project is about learning the Verilog-AMS programming language. It only makes sense to Verilog-AMS the official language for this project. It is getting its own project language file, starting here.");
      $finish;
    end
endmodule

// File info
// File type: Verilog-AMS source file (*.v *.vh)
// File version: 1 (2022, Sunday, November 6th at 11:34 pm PST)
// Line count (including blank lines and compiler line): 25

// End of script */
