// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 1
// For: seanpm2001/Learn-SystemVerilog
// About:
// I decided to make SystemVerilog the main project language file for this project (Seanpm2001/Learn-SystemVerilog) as SystemVerilog is the language this project is dedicated to, because this project is about learning the SystemVerilog programming language. It only makes sense to SystemVerilog the official language for this project. It is getting its own project language file, starting here.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 01'00000000 // Random data to test syntax
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: SystemVerilog source file (*.sv *.svh)
// File version: 1 (2022, Friday, September 23rd at 9:32 pm PST)
// Line count (including blank lines and compiler line): 16
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script
