// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 1
// For: Metro Techno / Traffic Light
// I decided to make Verilog the first project language file for this project (Seanpm2001/MetroTechno_Traffic) as Verilog is the primary language used for system programming on traffic lights running MetroTechno. C is used as a secondary laguage. Verilog comes first. It is getting its own project language file, starting here.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 01'00000000 // Random data to test syntax (also: 0 in binary)
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: Verilog source file (*.v *.vh)
// File version: 1 (2022, Wednesday, September 7th at 7:23 pm PST)
// Line count (including blank lines and compiler line): 15
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script
