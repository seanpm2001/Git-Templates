// Start of script */

// Project language file 1
// For: seanpm2001/Learn-Verilog
// About:
// I decided to make Verilog the main project language file for this project (Seanpm2001/Learn-Verilog) as Verilog is the language this project is dedicated to, because this project is about learning the Verilog programming language. It only makes sense to Verilog the official language for this project. It is getting its own project language file, starting here.

module main;
  initial
    begin
      $display("Project language file 1");
      $display("For: seanpm2001/Learn-Verilog");
      $display("About:");
      $display("I decided to make Verilog the main project language file for this project (Seanpm2001/Learn-Verilog) as Verilog is the language this project is dedicated to, because this project is about learning the Verilog programming language. It only makes sense to Verilog the official language for this project. It is getting its own project language file, starting here.");
      $finish;
    end
endmodule

// File info
// File type: Verilog source file (*.v *.vh)
// File version: 1 (2022, Saturday, November 5th at 10:52 pm PST)
// Line count (including blank lines and compiler line): 25

// End of script */
