// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 1
// For: SNU/2D/ProgrammingTools/IDE/SystemVerilog
// About:
// I decided to make SystemVerilog the main project language file for this project (SNU / 2D / Programming Tools / IDE / SystemVerilog) as this is a SystemVerilog IDE, and it needs its main language to be represented here.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 01'00000000 // Random data to test syntax
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: SystemVerilog source file (*.sv *.svh)
// File version: 1 (2022, Friday, September 23rd at 9:37 pm PST)
// Line count (including blank lines and compiler line): 16
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script
