// Start of script
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project language 40
// For: WacOS
// I decided to make SystemVerilog the fourtieth project language file for this project (Seanpm2001/WacOS) as SystemVerilog is a good language for machine instructions at direct programmable hardware level (such as FPGA devices) it can be used for some portions of this project. It is being included for software diversity reasons, and will be used for some portions of the project. It is getting its own project language file, starting here.
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`define PROJECT_LANG 40'00000100 // Random data to test syntax
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// File info:
// File type: SystemVerilog source file (*.sv *.svh)
// File version: 1 (Friday, 2021 December 24th at 4:31 pm)
// Line count (including blank lines and compiler line): 15
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// End of script

